// Twiddle factors for NTT
`define TWIDDLE_0 1
`define TWIDDLE_1 4150
`define TWIDDLE_2  1 // Continue defining all twiddle factors up to TWIDDLE_127
// ...
`define TWIDDLE_127  // Last twiddle factor